Your Hand Drawn Circuit's Netlist

V0 2 0 AC 45
D0 0 3 D1N4148
L0 1 3 45mH
R0 2 1 45

.tran 0.1ms 10ms
